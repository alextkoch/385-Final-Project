module graphics ( input logic [7:0] addr,
						output logic [31:0] data);

parameter[0:255][31:0] ROM = {

// tank up
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b11110000000000111100000000001111,
32'b11110000000000111100000000001111,
32'b10010000000000111100000000001001,
32'b10010000000000111100000000001001,
32'b11110000000000111100000000001111,
32'b11110000000000111100000000001111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11110000000000000000000000001111,
32'b11110000000000000000000000001111,

//tank left
32'b00001111111111111111111111111111,
32'b00001100110011001100110011001111,
32'b00001100110011001100110011001111,
32'b00001111111111111111111111111111,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b11111111111111111111111111111100,
32'b11111111111111111111111111111100,
32'b11111111111111111111111111111100,
32'b11111111111111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00000000001111111111111111111100,
32'b00001111111111111111111111111111,
32'b00001100110011001100110011001111,
32'b00001100110011001100110011001111,
32'b00001111111111111111111111111111,

//tank down
32'b11110000000000000000000000001111,
32'b11110000000000000000000000001111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b10011111111111111111111111111001,
32'b10011111111111111111111111111001,
32'b11110000000000111100000000001111,
32'b11110000000000111100000000001111,
32'b10010000000000111100000000001001,
32'b10010000000000111100000000001001,
32'b11110000000000111100000000001111,
32'b11110000000000111100000000001111,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,

//tank right
32'b11111111111111111111111111110000,
32'b11110011001100110011001100110000,
32'b11110011001100110011001100110000,
32'b11111111111111111111111111110000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111111111111111,
32'b00111111111111111111111111111111,
32'b00111111111111111111111111111111,
32'b00111111111111111111111111111111,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b00111111111111111111110000000000,
32'b11111111111111111111111111110000,
32'b11110011001100110011001100110000,
32'b11110011001100110011001100110000,
32'b11111111111111111111111111110000,

// bullet
32'b00000000000000000000000000000000, 
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000111100000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,

// brick
32'b11111111000011111110000011111111, 
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b00000000000000000000000000000000,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,
32'b11111111000011111110000011111111,

// bush; 0 is dark green, 1 is light green
32'b00000000000000000000000001110000,
32'b00000000000000000000000001110000,
32'b00000000000000000000000001110000,
32'b00000000110000000000000000000000,
32'b00000000110000000000000000000000,
32'b00000000110000000000000000000000,
32'b00001111111111111111111111111111,
32'b00001111111111111111111111111111,
32'b00001111111111111111111111111111,
32'b00001111111111111111111111111111,
32'b00001111111111110111111111111111,
32'b00001111111111110111111111111111,
32'b00001111111111110111110000011111,
32'b00001111111111110111110000011111,
32'b00001111111111110111110000011111,
32'b00111100111111111111111111111111,
32'b00111100111111111111111111111111,
32'b00111100111111111111111111111111,
32'b00111100111111111111111111111111,
32'b00001111111111111111111111110001,
32'b00001111111111111111111111111111,
32'b00001111111111111111111111111111,
32'b00001111111111111111111111111111,
32'b00001111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111110011111111111111111,
32'b00001111111110011111111111111111,
32'b00001111111110011111111111111111,
32'b00001111111110000000111111111111,

// Rock; 0 is darg gray, 1 is light gray
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11100000000000000000000000001100,
32'b11101111111111111111111111101100,
32'b11101111111111111111111111101100,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11101111111111111111111111100000,
32'b11100000000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11111100000000000000000000000000,
32'b11100000000000000000000000000000,
32'b11100000000000000000000000000000,


	};
	
	assign data = ROM[addr];

endmodule 
